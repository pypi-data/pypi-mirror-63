* test
v1 1 0 sin 0.5 0.5 4e9
r1 1 2 1
r2 2 0 1
.tran 0.1n 1n
.probe tran v(1) v(2) i(v1)
.option probe post=1
.end
