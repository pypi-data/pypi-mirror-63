* test
v1 1 0 DC 0.5 AC 1
r1 1 2 1
r2 2 0 1
c1 2 0 10p
.ac dec 20 1 1G
.probe ac v(1) v(2) i(v1)
.option probe post=1
.end
